/*
1.constraint restrict the random data generation to meaning values.
2.constraint are declarative and bidirectional code
syntax- constraint_identifier{constraiint expression[];}
*/
