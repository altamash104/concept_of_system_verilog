/*
1.It is a memory whose size is not known during compilation ,but instead is defined and expanded in as needed during the runtime.
2.A dynamic array is easily recognized by its empty square bracket[].
3.It is used in for small memory size upto range 1K to 1MB.
4.     declaration : bit [3:0] da[];
                      integer da[];
       memory allocation: da=new[4];
       da initializing :da={0,1,2,3} or '{0,1,2,3}
       dynamic array method: new[] Allocate the memory
       Return the size of an array : size()
       Delete all the elements of an array : delete()
       
*/

